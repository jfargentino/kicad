.title B&K 8103 hydrophone and its wire models
********************************************************************************
* 3.7nF 2.5GOhm with wire
* sensitivity -211dB 1V/uPa <-> 29uV/Pa <-> 0.1pC/Pa
*
* TODO simulate it and check C/R values for resonance freq and/or band pass
*      maybe a circuit topology could explain rx/tx assymetry ?
* 
* TODO a projector version, does it works to excit it and record in low
*      voltage to trace its bode ?
*
********************************************************************************
* Voltage source modelization
********************************************************************************
.subckt BK8103_V 1 2

* signal due to the ceramic deformation
* for a SPL of 60dB(1uPa), given the sensitivity, we should have 29nV
V1 4 2 DC 0 AC 30nV

* Equivalent capacitor of the ceramic
* given by C=Q/V and sensibility: 0.1pC/29uV = 3.448nF
C1 4 3 3.5nF

* Leakage resistor of the ceramic
R1 4 3 2.5G

* Equivalent resistance of the wire
R2 3 1 100m

* Equivalent capacitor of the wire
* Given by datasheet value less C1
C2 2 1 200pF

.ends BK8103_V

********************************************************************************
* Charge source modelization, BK8103_V Norton equivalent
********************************************************************************
.subckt BK8103_I 1 2

* TODO Norton equivalent of V1
I1 2 3 DC 0 AC 100pA
C1 2 3 3.5nF
R1 2 3 2.5G
R2 3 1 100m
C2 2 1 200pF

.ends BK8103_I

********************************************************************************
* Transducer+wire modelization, passive
********************************************************************************
.subckt BK8103_P 1 2

C1 2 3 3.5nF
R1 2 3 2.5G
R2 3 1 100m
C2 2 1 200pF

.ends BK8103_P

********************************************************************************
* Just sources useful for some simulations
********************************************************************************
.subckt BK8103_SIMU_V 1 2
V1 1 2 DC 0u AC 1u
.ends BK8103_SIMU_V

.subckt BK8103_SIMU_I 1 2
I1 1 2 DC 0u AC 1u
.ends BK8103_SIMU_I

********************************************************************************
