.title B&K 8103 hydrophone and its wire models
********************************************************************************
* 3.7nF 2.5GOhm with wire
* sensitivity -211dB 1V/uPa <-> 29uV/Pa <-> 0.1pC/Pa
*
* TODO simulate it and check C/R values for resonance freq and/or band pass
*      maybe a circuit topology could explain rx/tx assymetry ?
********************************************************************************
* Charge source modelization
********************************************************************************
.subckt BK8103_Q 1 2

* signal due to the ceramic deformation
* TODO transpose 0.1pC/Pa into a realistic current (i = dq/dt)
I1 2 3 DC 0 AC 100pA

* Equivalent capacitor of the ceramic
* given by C=Q/V and sensibility: 0.1pC/29uV = 3.448nF
C1 2 3 3.5nF

* Leakage resistor for the ceramic
R1 2 3 2.5G

* Equivalent resistance of the wire
R2 3 1 100m

* Equivalent capacitor of the wire
* Given by datasheet value less C1
C2 2 1 200pF

.ends BK8103_Q

********************************************************************************
* Voltage source modelization
********************************************************************************
.subckt BK8103_V 1 2

* signal due to the ceramic deformation
* for a SPL of 60dB(1uPa),  given the sensitivity, we should have 29nV
V1 4 2 DC 0 AC 30nV

* Equivalent capacitor of the ceramic
* given by C=Q/V and sensibility: 0.1pC/29uV = 3.448nF
C1 4 3 3.5nF

* Leakage resistor for the ceramic
R1 4 3 2.5G

* Equivalent resistance of the wire
R2 3 1 100m

* Equivalent capacitor of the wire
* Given by datasheet value less C1
C2 2 1 200pF

.ends BK8103_V
********************************************************************************

