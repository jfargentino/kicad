* OPA132 PSpice Model (PSpice format)
********************************************
**  This file was created by TINA        **
**    (c) 1996-2006 DesignSoft, Inc.   **
********************************************
* OPA132 REV A  CREATED BY MAREK LIS
* GREEN-LIS MACRO-MODEL ARCHITECTURE
* DECEMBER 20, 2013
*
* THIS MACROMODEL HAS BEEN OPTIMIZED TO MODEL THE AC, DC, NOISE, AND TRANSIENT RESPONSE PERFORMANCE WITHIN
* THE DEVICE DATA SHEET SPECIFIED LIMITS. CORRECT OPERATION OF THIS MACROMODEL HAS BEEN VERIFIED ON DESIGNSOFT
* TINA VERSION 7.0.80.224 SF. FOR HELP WITH OTHER ANALOG SIMULATION SOFTWARE, PLEASE CONSULT THE SOFTWARE SUPPLIER.
*
* COPYRIGHT 2011 BY TEXAS INSTRUMENTS CORPORATION
*
* BEGIN MODEL OPA132
*
*GREEN-LIS MACRO-MODEL SIMULATED TYPICAL PARAMETERS:
*
*OPEN LOOP GAIN AND PHASE VS FREQUENCY WITH RL AND CL EFFECTS
*INPUT COMMON MODE REJECTION WITH FREQUENCY
*POWER SUPPLY REJECTION WITH FREQUENCY
*INPUT IMPEDANCE VS FREQUENCY
*OUTPUT IMPEDANCE VS FREQUENCY AND OUTPUT CURRENT
*INPUT VOLTAGE NOISE VS FREQUENCY
*INPUT CURRENT NOISE VS FREQUENCY
*OUTPUT VOLTAGE SWING VS OUTPUT CURRENT
*SHORT-CIRCUIT OUTPUT CURRENT
*QUIESCENT CURRENT VS SUPPLY VOLTAGE
*SETTLING TIME VS CAPACITIVE LOAD
*SLEW RATE
*SMALL SIGNAL OVERSHOOT VS CAPACITIVE LOAD
*LARGE SIGNAL RESPONSE
*OVERLOAD RECOVERY TIME
*INPUT BIAS CURRENT
*INPUT VOLTAGE OFFSET
*INPUT COMMON MODE RANGE
*OUTPUT CURRENT COMING THROUGH THE SUPPLY RAILS

.SUBCKT OPA132 +IN -IN V+ V- Vout
V7          15 56 2.8
Vos         28 47 -100.1U
V11         58 59 100M
V10         60 61 100M
V6          11 66 10
V5          67 11 10
V4          63 65 10
V1          64 62 10
V9          78 16 2.8
IS2         V+ 28 5P
IS1         V+ V- 4M
IS3         52 V- -7P
V3          82 11 40
V2          11 83 47
R37         29 30 100MEG
C4          31 29  1.00000000000000E-0016 IC=0
C1          11 32 1N IC=0
EVCVS1      10 11 7 33  -1
R38         32 34 10
VCCVS2_in   33 8
HCCVS2      34 11 VCCVS2_in   1K
XU7         32 11 33 30 VC_RES_0
C25         10 31 2P IC=0
C24         10 9 90N IC=0
R32         9 31 10.5K
R31         31 30 100MEG
R30         10 31 500K
EVCVS2      30 11 11 31  20MEG
SW14        9 10 12 11  S_VSWITCH_1
SW13        10 9 11 13  S_VSWITCH_2
XR105       14 11 RNOISE_FREE_0
XR105_2     35 11 RNOISE_FREE_1
R24         11 20 1K
R17         11 21 1K
R11         11 36 1K
R10         11 37 1K
R9          11 12 1K
R8          11 13 1K
L4          11 38 17M IC=0
L1          39 11 1F IC=0
R2          39 40 1
GVCCS8      11 40 11 41  1
XR109       42 11 RNOISE_FREE_1
C3          42 11 3F IC=0
GVCCS4      11 42 25 11  1U
C2          43 11 3F IC=0
XR109_2     43 11 RNOISE_FREE_2
GVCCS3      11 43 42 11  1M
R4          44 23 10M
CinDiff     45 46 2P IC=0
CinpCM      46 11 5P IC=0
CinnCM      11 45 5P IC=0
XIn11       47 45 FEMT_0
L2          48 11 1F IC=0
XR109_3     25 11 RNOISE_FREE_1
XR109_4     49 11 RNOISE_FREE_1
XVn11       46 47 VNSE_0
XU14        50 11 51 52 VCVS_LIMIT_0
L3          53 11 350U IC=0
R1          48 50 1
GVCCS2      11 50 11 54  1
XU13        15 55 IDEAL_D_0
EVCVS5      56 11 V- 11  1
C11         49 11 4F IC=0
XR109_5     24 11 RNOISE_FREE_2
GVCCS12     11 25 49 11  1U
XU5         17 11 V+ 18 VCVS_LIMIT_1
XU6         11 17 19 V- VCVS_LIMIT_2
C15         V+ V- 10P IC=0
C22         11 22 1P IC=0
R29         22 14 1
C23         11 26 1P IC=0
C9          57 11 10P IC=0
R26         57 17 10
C21         11 12 1P IC=0
C20         11 13 1P IC=0
C19         20 11 1P IC=0
C17         21 11 1P IC=0
C16         11 36 1P IC=0
C12         37 11 1P IC=0
R13         7 26 1
R36         26 61 1M
R35         26 59 1M
SW12        62 58 20 11  S_VSWITCH_3
SW11        60 63 11 21  S_VSWITCH_4
R34         26 64 1K
R33         26 65 1K
SW10        67 14 22 11  S_VSWITCH_5
SW9         14 66 11 22  S_VSWITCH_6
R25         68 20 1
R19         69 21 1
R16         70 36 1
R14         71 37 1
R12         72 12 1
R7          73 13 1
R5          74 24 10M
R6          75 14 10M
R15         0 11 100MEG
C13         24 11 1F IC=0
GVCCS1      11 24 43 11  1M
GIsinking   V- 11 76 11  1M
GIsourcing  V+ 11 77 11  1M
R23         76 11 10K
SW7         17 76 57 11  S_VSWITCH_7
R21         11 77 10K
SW8         17 77 57 11  S_VSWITCH_8
SW4         75 72 12 11  S_VSWITCH_9
SW3         73 75 11 13  S_VSWITCH_10
XU3         63 27 73 11 VCVS_LIMIT_3
XU1         62 27 72 11 VCVS_LIMIT_3
SW2         44 68 20 11  S_VSWITCH_11
SW1         69 44 11 21  S_VSWITCH_12
XU8         28 V+ IDEAL_D_1
XU12        V- 28 IDEAL_D_1
EVCVS6      78 11 V+ 11  1
R22         79 55 100
EVCVS4      79 11 28 11  1
XU2         55 16 IDEAL_D_0
SW6         74 70 36 11  S_VSWITCH_13
SW5         71 74 11 37  S_VSWITCH_14
XU26        55 52 11 80 VCCS_LIMIT_0
XU4         80 11 11 14 VCCS_LIMIT_1
LPSR        81 11 3.16M IC=0
XVCVSPSRR   40 11 51 45 VCVS_LIMIT_4
XU22        82 17 69 11 VCVS_LIMIT_5
XU21        83 17 68 11 VCVS_LIMIT_5
XU20        19 Vout 70 11 VCVS_LIMIT_5
XU19        18 Vout 71 11 VCVS_LIMIT_6
XU11        V- 52 IDEAL_D_1
XU10        52 V+ IDEAL_D_1
C10         23 11 1F IC=0
C5          25 11 4F IC=0
XR109_6     23 11 RNOISE_FREE_2
GVCCS15     11 23 24 11  1M
GVCCS10     11 49 35 11  1U
R20         +IN 46 100
R18         -IN 45 100
GVCCS6      11 35 27 11  1U
XR102       84 85 RNOISE_FREE_1
XR101       86 84 RNOISE_FREE_1
C6          84 0 1 IC=0
XR105_3     27 11 RNOISE_FREE_1
XR103       11 80 RNOISE_FREE_1
EVCVS34     11 0 84 0  1
RPSR        81 41 1
GVCCS11     11 41 V+ V-  5U
RCM         53 54 1
EVCVS29     86 0 V+ 0  1
EVCVS28     85 0 V- 0  1
GVCCS7      11 54 28 11  10U
VCCVS1_in   8 Vout
HCCVS1      17 11 VCCVS1_in   1K
GVCCS5      11 27 14 11  1U
Ccc         14 11 3.8U IC=0
EVCVS3      7 11 23 11  1
.MODEL S_VSWITCH_1 VSWITCH (RON=1 ROFF=100MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_2 VSWITCH (RON=1 ROFF=100MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_3 VSWITCH (RON=1 ROFF=10MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_4 VSWITCH (RON=1 ROFF=10MEG VON=100M VOFF=-100M)
.MODEL S_VSWITCH_5 VSWITCH (RON=10M ROFF=100MEG VON=150 VOFF=130)
.MODEL S_VSWITCH_6 VSWITCH (RON=10M ROFF=100MEG VON=150 VOFF=130)
.MODEL S_VSWITCH_7 VSWITCH (RON=1M ROFF=10MEG VON=-10M VOFF=0)
.MODEL S_VSWITCH_8 VSWITCH (RON=1M ROFF=10MEG VON=10M VOFF=0)
.MODEL S_VSWITCH_9 VSWITCH (RON=1 ROFF=10MEG VON=1 VOFF=-1)
.MODEL S_VSWITCH_10 VSWITCH (RON=1 ROFF=10MEG VON=1 VOFF=-1)
.MODEL S_VSWITCH_11 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_12 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_13 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.MODEL S_VSWITCH_14 VSWITCH (RON=1 ROFF=1G VON=10 VOFF=-10)
.ENDS


*VOLTAGE CONTROLLED RESISTOR
.SUBCKT VC_RES_0  1      2      3    4
*              VC+    VC-   RES1 RES2
ERES 3 40 VALUE = {(I(VSENSE) * (ABS(V(1,2))*ABS(V(1,2))*0.000352-0.02359*ABS(V(1,2))+0.5922))*140000*24200*50*2/414500}
VSENSE 40 4 DC 0
.ENDS VC_RES_0


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_0  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E4
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_0


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_1  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E6
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_1


* NOISELESS RESISTOR
.SUBCKT RNOISE_FREE_2  1 2
*ROHMS = VALUE IN OHMS OF NOISELESS RESISTOR
.PARAM ROHMS=1E3
ERES 1 3 VALUE = { I(VSENSE) * ROHMS }
RDUMMY 30 3 1
VSENSE 30 2 DC 0V
.ENDS RNOISE_FREE_2


* BEGIN PROG NSE FEMTO AMP/RT-HZ
.SUBCKT FEMT_0  1 2
* BEGIN SETUP OF NOISE GEN - FEMPTOAMPS/RT-HZ
* INPUT THREE VARIABLES
* SET UP INSE 1/F
* FA/RHZ AT 1/F FREQ
.PARAM NLFF=.001
* FREQ FOR 1/F VAL
.PARAM FLWF=0.001
* SET UP INSE FB
* FA/RHZ FLATBAND
.PARAM NVRF=0.1
* END USER INPUT
* START CALC VALS
.PARAM GLFF={PWR(FLWF,0.25)*NLFF/1164}
.PARAM RNVF={1.184*PWR(NVRF,2)}
.MODEL DVNF D KF={PWR(FLWF,0.5)/1E11} IS=1.0E-16
* END CALC VALS
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVNF
D2 8 0 DVNF
E1 3 6 7 8 {GLFF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNVF}
R5 5 0 {RNVF}
R6 3 4 1E9
R7 4 0 1E9
G1 1 2 3 4 1E-6
C1 1 0 1E-15
C2 2 0 1E-15
C3 1 2 1E-15
.ENDS
* END PROG NSE FEMTO AMP/RT-HZ


* BEGIN PROG NSE NANO VOLT/RT-HZ
.SUBCKT VNSE_0  1 2
* BEGIN SETUP OF NOISE GEN - NANOVOLT/RT-HZ
* INPUT THREE VARIABLES
* SET UP VNSE 1/F
* NV/RHZ AT 1/F FREQ
.PARAM NLF=83
* FREQ FOR 1/F VAL
.PARAM FLW=1
* SET UP VNSE FB
* NV/RHZ FLATBAND
.PARAM NVR=7.5
* END USER INPUT
* START CALC VALS
.PARAM GLF={PWR(FLW,0.25)*NLF/1164}
.PARAM RNV={1.184*PWR(NVR,2)}
.MODEL DVN D KF={PWR(FLW,0.5)/1E11} IS=1.0E-16
* END CALC VALS
I1 0 7 10E-3
I2 0 8 10E-3
D1 7 0 DVN
D2 8 0 DVN
E1 3 6 7 8 {GLF}
R1 3 0 1E9
R2 3 0 1E9
R3 3 6 1E9
E2 6 4 5 0 10
R4 5 0 {RNV}
R5 5 0 {RNV}
R6 3 4 1E9
R7 4 0 1E9
E3 1 2 3 4 1
C1 1 0 1E-15
C2 2 0 1E-15
C3 1 2 1E-15
.ENDS
* END PROG NSE NANOV/RT-HZ


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_0  VC+ VC- VOUT+ VOUT-
*             
.PARAM GAIN = 1
.PARAM VPOS = 10M
.PARAM VNEG = -10M
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS VCVS_LIMIT_0


*TG IDEAL DIODE
.SUBCKT IDEAL_D_0  A C
D1 A C DNOM
.MODEL DNOM D (TT=10P CJO=1E-18 IS=1E-15 RS=1E-3)
.ENDS IDEAL_D_0


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_1  VC+ VC- VOUT+ VOUT-
*             

E1 VOUT+ VOUT- TABLE {ABS(V(VC+,VC-))} = (0.0,0.9)(20,2.0)(30,2.6)(39.9,3.7)
.ENDS VCVS_LIMIT_1



*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_2  VC+ VC- VOUT+ VOUT-
*             

E1 VOUT+ VOUT- TABLE {ABS(V(VC+,VC-))} = (0.0,0.3)(3,0.3)(5,0.5)(6,0.9)(46.9,3.3)
.ENDS VCVS_LIMIT_2


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_3  VC+ VC- VOUT+ VOUT-
*             
.PARAM GAIN = 100
.PARAM VPOS = 6000
.PARAM VNEG = -6000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS VCVS_LIMIT_3


*TG IDEAL DIODE
.SUBCKT IDEAL_D_1  A C
D1 A C DNOM
.MODEL DNOM D (TT=10P CJO=1E-18 IS=1E-15 RS=1E-3)
.ENDS IDEAL_D_1


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_0  VC+ VC- IOUT+ IOUT-
*             
.PARAM GAIN = 1M
.PARAM IPOS = .5
.PARAM INEG = -.5
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS VCCS_LIMIT_0


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCCS_LIMIT_1  VC+ VC- IOUT+ IOUT-
*             
.PARAM GAIN = 200M
.PARAM IPOS = 76
.PARAM INEG = -76
G1 IOUT+ IOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),INEG,IPOS)}
.ENDS VCCS_LIMIT_1


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_4  VC+ VC- VOUT+ VOUT-
*             
.PARAM GAIN = -1
.PARAM VPOS = 10M
.PARAM VNEG = -10M
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS VCVS_LIMIT_4


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_5  VC+ VC- VOUT+ VOUT-
*             
.PARAM GAIN = 100
.PARAM VPOS = 5000
.PARAM VNEG = -5000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS VCVS_LIMIT_5


*VOLTAGE CONTROLLED SOURCE WITH LIMITS
.SUBCKT VCVS_LIMIT_6  VC+ VC- VOUT+ VOUT-
*            
.PARAM GAIN = 100
.PARAM VPOS = 5000
.PARAM VNEG = -5000
E1 VOUT+ VOUT- VALUE={LIMIT(GAIN*V(VC+,VC-),VNEG,VPOS)}
.ENDS VCVS_LIMIT_6

.END
