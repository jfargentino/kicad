.title B&K 8103 hydrophone and its wire model
********************************************************************************
.subckt BK8103 1 2

* signal due to the ceramic deformation
Isignal 2 4 AC 100p

* Equivalent capacitor of the ceramic
Chydro 3 4 3.2n

* Leakage resistor for the ceramic
Rhydro 3 2 2.5G

* Equivalent capacitor of the wire
Cwire 3 2 500p

* Equivalent resistance of the wire
Rwire 1 3 100m

********************************************************************************
.ends BK8103

